----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:50:23 03/26/2018 
-- Design Name: 
-- Module Name:    I2C - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------



---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY I2C IS 
	PORT (RESET 		: IN 	STD_LOGIC;
			CLK_2M		: IN	STD_LOGIC;
		  SCL, SDATA_DIR: OUT 	STD_LOGIC;
			SDATA 		: INOUT STD_LOGIC);
END I2C;

ARCHITECTURE Behavioral OF I2C IS
SIGNAL REGISTER_CHANGED			: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL INSTRUCTION_CHANGED	 	: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL DATA_CHANGED				: STD_LOGIC_VECTOR (7 DOWNTO 0); 
SIGNAL DATA_REALWRITE			: STD_LOGIC_VECTOR (7 DOWNTO 0); 
SIGNAL COUNT					: INTEGER RANGE 0 TO 9;
SIGNAL COUNT_CONTROL			: INTEGER RANGE 0 TO 63;
SIGNAL COUNT_ACK				: INTEGER RANGE 0 TO 3;
SIGNAL COUNT_DATAWRITED			: INTEGER RANGE 0 TO 3;
SIGNAL COUNT_10HZ				: INTEGER RANGE 0 TO 204799;
SIGNAL CLK_10HZ 				: STD_LOGIC;
SIGNAL CLK_200K					: STD_LOGIC;
SIGNAL CLK_100K 				: STD_LOGIC;
SIGNAL CLK_50K 					: STD_LOGIC;

TYPE STATETYPE IS (NORMAL_STATE, WAITACK_STATE, WRITEDATA_STATE, END_STATE);
SIGNAL I2CCONTROLSTATE 		: STATETYPE;
BEGIN
REGISTER_CHANGED		<="01010000";
INSTRUCTION_CHANGED		<="10100100";
DATA_CHANGED			<="00111000";

PROCESS(CLK_2M) --从2M时钟产生200K,100K和50K时钟信号
BEGIN
	IF (CLK_2M'EVENT AND CLK_2M='1') THEN
		IF(COUNT_10HZ=204799) THEN COUNT_10HZ<=0;
			CLK_10HZ <= NOT CLK_10HZ;
		ELSE COUNT_10HZ <=COUNT_10HZ+1;
		END IF;
	END IF;
END PROCESS;


PROCESS(CLK_2M,RESET) 
BEGIN
	IF (RESET='1') THEN COUNT <=0;CLK_200K<='0';
	  ELSIF (CLK_2M'EVENT AND CLK_2M='1') THEN
	  	IF(COUNT=9) THEN COUNT<=0; CLK_200K<= NOT CLK_200K;
	  		ELSE COUNT<=COUNT +1;
		END IF;
	END IF;
END PROCESS;

PROCESS(CLK_200K,RESET) 
BEGIN
	IF (RESET='1') THEN CLK_100K<='0';
	  ELSIF (CLK_200K'EVENT AND CLK_200K='1') THEN
	  	    CLK_100K<= NOT CLK_100K;
	END IF;
END PROCESS;
 
PROCESS(CLK_100K,RESET) 
BEGIN
	IF (RESET='1') THEN CLK_50K<='0';
	  ELSIF (CLK_100K'EVENT AND CLK_100K='1') THEN
	  	    CLK_50K<= NOT CLK_50K;
	END IF;
END PROCESS;
SCL<=CLK_50K;


PROCESS (RESET,CLK_200K)--产生写 WR 寄存器的时序
BEGIN
	IF(RESET='1')
		THEN COUNT_CONTROL<=0;
	ELSIF (CLK_200K'EVENT AND CLK_200K= '1') THEN
	 CASE I2CCONTROLSTATE IS
		WHEN NORMAL_STATE	=>	COUNT_CONTROL<=COUNT_CONTROL +1 ;
		WHEN WAITACK_STATE 	=>	COUNT_CONTROL<= 0;
		WHEN WRITEDATA_STATE=>	COUNT_CONTROL<=COUNT_CONTROL +1 ;
		WHEN END_STATE 		=>	COUNT_CONTROL<=	0;
		WHEN OTHERS 		=> 	NULL;
	 END CASE;
	END IF;
END PROCESS ;

PROCESS (RESET,CLK_200K)
BEGIN
	IF(RESET='1') THEN SDATA<='1' ;SDATA_DIR<='1';
		I2CCONTROLSTATE <= NORMAL_STATE;
	ELSIF(CLK_200K'EVENT AND CLK_200K='0') THEN
	CASE I2CCONTROLSTATE IS
	 WHEN NORMAL_STATE =>
		IF(COUNT_CONTROL=1) THEN SDATA <='0';
			ELSIF(COUNT_CONTROL=3) THEN
				SDATA<=REGISTER_CHANGED(7);
			ELSIF(COUNT_CONTROL=7) THEN
				SDATA<=REGISTER_CHANGED(6);
			ELSIF (COUNT_CONTROL=11) THEN
				SDATA<=REGISTER_CHANGED(5);
			ELSIF (COUNT_CONTROL=15) THEN
				SDATA<=REGISTER_CHANGED(4);
			ELSIF (COUNT_CONTROL=19) THEN
				SDATA<=REGISTER_CHANGED(3);
			ELSIF (COUNT_CONTROL=23) THEN
				SDATA<=REGISTER_CHANGED(2) ;
			ELSIF (COUNT_CONTROL=27) THEN
				SDATA<=REGISTER_CHANGED(1) ;
			ELSIF (COUNT_CONTROL=31) THEN
				SDATA<=REGISTER_CHANGED(0) ;
			ELSIF (COUNT_CONTROL=35) THEN
				SDATA<='Z';
				I2CCONTROLSTATE<=WAITACK_STATE;
		END IF;
			SDATA_DIR <='1';
	 WHEN WAITACK_STATE =>
			SDATA_DIR <='0';SDATA<='Z';
		IF (SDATA='0') THEN COUNT_ACK <=COUNT_ACK +1;
		END IF;
		IF (COUNT_ACK=2) THEN 
			IF (COUNT_DATAWRITED=0) THEN 
				I2CCONTROLSTATE <=	WRITEDATA_STATE;
				DATA_REALWRITE	<=	INSTRUCTION_CHANGED;
				COUNT_DATAWRITED<=	COUNT_DATAWRITED +1;
			ELSIF (COUNT_DATAWRITED=1) THEN
				I2CCONTROLSTATE <=	WRITEDATA_STATE;
				DATA_REALWRITE	<=	DATA_CHANGED;
				COUNT_DATAWRITED<=	COUNT_DATAWRITED +1;
			ELSIF (COUNT_DATAWRITED=2) THEN 
				COUNT_DATAWRITED<=	0;
				I2CCONTROLSTATE <=	END_STATE;
			END IF;
		ELSE I2CCONTROLSTATE <= WAITACK_STATE;
		END IF;
	 WHEN WRITEDATA_STATE =>
				IF(COUNT_CONTROL=1) THEN
					SDATA<=DATA_REALWRITE (7) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=5) THEN
					SDATA<=DATA_REALWRITE (6) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=9) THEN
					SDATA<=DATA_REALWRITE (5) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=13) THEN
					SDATA<=DATA_REALWRITE (4) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=17) THEN
					SDATA<=DATA_REALWRITE (3) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=21) THEN
					SDATA<=DATA_REALWRITE (2) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=25) THEN
					SDATA<=DATA_REALWRITE (1) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=29) THEN
					SDATA<=DATA_REALWRITE (0) ;
					SDATA_DIR<='1';
				ELSIF(COUNT_CONTROL=33) THEN
					SDATA<='Z';
					I2CCONTROLSTATE<=WAITACK_STATE;
					COUNT_ACK<=0;
					SDATA_DIR<='0';
				END IF;
	 WHEN END_STATE=>SDATA<='1';
					SDATA_DIR<='1';
	 WHEN OTHERS =>NULL;
	END CASE;
	END IF;
END PROCESS;
END Behavioral; 









